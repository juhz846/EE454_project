module Conv2d #(
    parameter window_size,
    parameter channels,
    parameter neurons
) (
    
    
);
    
endmodule


module MaxPool #(
    parameters
) (
    ports
);
    
endmodule

module FC #(
    parameters
) (
    ports
);
    
endmodule


module CNN #(
    parameters
) (
    ports
);
    
endmodule